----------------------------------------------------------------------------------
-- Company:MPOR 
-- Engineer:maher and ashour
-- 
-- Create Date:    15:35:52 02/14/2019 
-- Design Name: 
-- Module Name:    ins_mem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_logic_unsigned.ALL;
use IEEE.STD_LOGIC_arith.ALL;
entity ins_mem is
generic(data_width: integer:=32;
        add_bits: integer := 5);
    Port ( pc : in  STD_LOGIC_VECTOR ( add_bits-1 downto 0);
           instruction : out  STD_LOGIC_VECTOR (data_width-1 downto 0));
end ins_mem;



architecture Behavioral of ins_mem is

type ins_type is array (0 to 2047) of std_logic_vector(data_width-1 downto 0);

signal ins_mem : ins_type;

begin

ins_mem <= ("00000000000000000000010000000000",
"00000000010001000100010000000000",
"00000000110011001100010000000000",
"10000000000000000000000000000101",
"10000000010001000000000001100001",
"00000000000001001000000000000000",
"10000000110011000000000001100110",
"01000100000000000000000000001011",
"11000000010011000000000000000010",
"00000000000000000000010000000000",
"00111100000000000000000000000000",
"10110100000001000000000000000000",
"10110100000010000000000000000000",
"10111000000001000000000000000000",
"10111000000010000000000000000000",
"01001000000000000000000000000000",
"01000100000000000000000110101101",
"10010011111111000000000000000000",
"10000011111111000000000001011100",
"11000001101111000000000000000110",
"10000011111111000000000000000001",
"11000001101111000000000000000111",
"10000011111111000000000000000001",
"11000001101111000000000000001000",
"01000000000000000000000000000110",
"10010011111111000000000000000000",
"10000011110001000000000000000001",
"01000000000000000000000000011100",
"10010011111111000000000000000000",
"10000011110001000000000000000010",
"01000000000000000000000000011100",
"10010011111111000000000000000000",
"10000011110001000000000000000011",
"01000000000000000000000000011100",
"10010000100010000000000000000000",
"10110000000111000000000000000010",
"10110100000001000000000000000000",
"10010000010001000000000000000000",
"10000001110001000000000000000000",
"01000100000000000000001011010001",
"10111000000001000000000000000000",
"01000000000000000000000000110101",
"10010011111111000000000000000000",
"10010111111111000000000000000010",
"11000100011111000000000000000101",
"10000011111111000000000000000101",
"11000000111111000000000001100001",
"11000001000111000000000001101101",
"01000000000000000000000000110101",
"10010011111111000000000000000000",
"10010111111111000000000000000011",
"11000000111111000000000001011100",
"11000001000111000000000001101000",
"10010010001000000000000000000000",
"10010110001000000000000000000001",
"01000100000000000000000111010111",
"10010011111111000000000000000000",
"10000011111111000000000001011011",
"11000101101111000000000000001000",
"10010011111111000000000000000000",
"10010111111111000000000000000001",
"11000100011111111111111111111000",
"10000011111111000000000000000001",
"11000000101111111111111111110110",
"10000000100010000000000000000001",
"01000000000000000000000000110101",
"10010011001100000000000000000000",
"10010011111111000000000000000000",
"10010111111111000000000000000011",
"11000010001111000000000001000001",
"10010010011001000000000000000000",
"00000010000000111100000000000000",
"10000111111111000000000000000001",
"10110011111010000000000000000000",
"10000110001111000000000000000011",
"10110011110101000000000000001010",
"10010011111111000000000000000000",
"10010111111111000000000000000100",
"11000110011111000000000000000011",
"10000010001000000000000000000001",
"01000000000000000000000001000011",
"10110100001010000000000000000000",
"10010010101010000000000011111111",
"11000101101010000000000000101000",
"10010010111011000000000000000000",
"10010110111011000000000000000001",
"10010011111111000000000000000000",
"11000011111001000000000000000100",
"10100010111011000000000000000000",
"10000011111111000000000000000001",
"01000000000000000000000001010111",
"10110100000101000000000000000000",
"00000010110101010101000000000000",
"11000010110101000000000000011101",
"10111000000101000000000000000000",
"00000001011011010101010000000000",
"10010011111111000000000000000000",
"10000011111111000000000000001010",
"00000011111000111100000000000000",
"10000111111111000000000000000011",
"10101111110101000000000000000000",
"10000001000100000000000000000001",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10110100001000000000000000000000",
"10110100001010000000000000000000",
"10010011111111000000000000000000",
"10010111111111000000000000000001",
"11000110001111000000000000000101",
"10010010101010000000000000000000",
"10010110101010000000000000000011",
"00000010101001000100010000000000",
"01000000000000000000000001110100",
"10010010101010000000000000000000",
"10010110101010000000000000000111",
"00000010101001000100010000000000",
"10000001100000000000000000000000",
"01000100000000000000001010111001",
"10111000001010000000000000000000",
"10111000001000000000000000000000",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"10010111001100000000000000000001",
"10111000001010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10100110101010000000000000000000",
"10000010011001000000000000000001",
"01000000000000000000000001001100",
"10010011111111000000000000000000",
"10011011111111000000000000000001",
"11000011001111111111111110011011",
"10000000110011000000000000000001",
"10110100001111000000000000000000",
"10000000111111000000000000000000",
"01000100000000000000001010100101",
"10111000001111000000000000000000",
"01000000000000000000000000100011",
"01000100000000000000001001011100",
"01000100000000000000001011000101",
"10000011101110000000000000000001",
"10010011111111000000000000000000",
"10000011111111000000000000001010",
"10000111111111000000000000000001",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10101111110000000000000000000000",
"10000111111111000000000000000001",
"10101111110000000000000000000000",
"10111000000000000000000000000000",
"01000000000000000000000000000100",
"01000100000000000000001001000001",
"01000100000000000000001011000101",
"10000011101110000000000000000001",
"10010011111111000000000000000000",
"10000011111111000000000000001010",
"10000111111111000000000000000001",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10101111110000000000000000000000",
"10000111111111000000000000000001",
"10101111110000000000000000000000",
"10111000000000000000000000000000",
"01000000000000000000000000000100",
"00111100000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"11010000000000000000000000000000",
"01000100000000000000000101001010",
"10000000000000000000000000111000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000001100",
"01000100000000000000000100011111",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000110",
"01000100000000000000000100011111",
"10010000000000000000000000000000",
"10000000000000000000000001001000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001101",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000010001111",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"10010011111111000000000000000000",
"10000011111111000000000000001000",
"10110011110101000000000000000000",
"10010001010101000000000000001111",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000110111000000000000010011",
"11000000101111000000000000000100",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000100000011",
"10110000000110000000000000000000",
"10010000100010000000000000000000",
"10010100100010000000000011111111",
"10001000111010000000000000001000",
"10010011111111000000000000000000",
"11000011111010000000000000000100",
"10100101100110000000000000000000",
"10000110101010000000000000000001",
"01000000000000000000000100001111",
"00000000100110011001000000000000",
"10110100000001000000000000000000",
"10010000010001000000000000000000",
"00000000010110000101010000000000",
"01000100000000000000001011100100",
"10111000000001000000000000000000",
"10111000000101000000000000000000",
"10111000000001000000000000000000",
"10111000000010000000000000000000",
"10111000000011000000000000000000",
"10111000000110000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"11010000000000000000000000000000",
"10010100000000000000000100000000",
"11010000000000000000000000000000",
"01000100000000000000000100110011",
"10010000000000000000000011111111",
"11010000000000000000000000000000",
"01000100000000000000000100111110",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"11010000000000000000000000000000",
"10010100000000000000001100000000",
"11010000000000000000000000000000",
"01000100000000000000000100110011",
"10010000000000000000111011111111",
"11010000000000000000000000000000",
"01000100000000000000000100111110",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000000011001",
"10010000010001000000000000000000",
"11000000000001000000000000000011",
"10000100000000000000000000000001",
"01000000000000000000000100111000",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001100100",
"10010000010001000000000000000000",
"11000000000001000000000000000100",
"01000100000000000000000100110011",
"10000100000000000000000000000001",
"01000000000000000000000101000011",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000000010100",
"10010000010001000000000000000000",
"11000000010000000000000000000100",
"01000100000000000000000100111110",
"10000100000000000000000000000001",
"01000000000000000000000101001111",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000000001000",
"10010000010001000000000000000000",
"11000000010000000000000000000100",
"01000100000000000000000101001010",
"10000100000000000000000000000001",
"01000000000000000000000101011011",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000110001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000111010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000101",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001011001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000010010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000110010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000111010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001101",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000011010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000110011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000111010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000100",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000100000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000010010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000100000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000011010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000100000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000010000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10110100000011000000000000000000",
"10110100000100000000000000000000",
"10110100000101000000000000000000",
"10010000000000000000000000000000",
"11010000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"10010000010001000000000000000000",
"10000000010001000000000000111111",
"11000100000001111111111111111001",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000000000001111111111111111011",
"01000100000000000000000101010110",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000000000001111111111111110111",
"10010000000000000000000000000000",
"10000000000000000011110000000000",
"11010000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000100000001000000000000100101",
"10010000000000000000000000000000",
"10000000000000000101110000000000",
"11010000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000100000001000000000000011110",
"10010000000000000000000000000000",
"10000000000000000110110000000000",
"11010000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000100000001000000000000011000",
"10010000000000000000000000000000",
"10000000000000000111010000000000",
"11010000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000100000001000000000000010010",
"10010000000000000000000000000000",
"10000000000000000111100000000000",
"11010000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"10000000000000000000000000000000",
"00101100000000000000000000000000",
"10010000000000000000000000111111",
"11000100000001000000000000001100",
"10010000100010000000000000000000",
"01000000000000000000001000101011",
"10010000100010000000000000000000",
"10000000100010000000000000000110",
"01000000000000000000001000101011",
"10010000100010000000000000000000",
"10000000100010000000000000001100",
"01000000000000000000001000101011",
"10010000100010000000000000000000",
"10000000100010000000000000010010",
"01000000000000000000001000101011",
"10010000100010000000000000000000",
"10000000100010000000000000011000",
"10010000110011000000000000000000",
"10010001000100000000000000000000",
"10010001010101000000000000000000",
"10000000110011000000000000000001",
"10110100000000000000000000000000",
"00000000000011000001000000000000",
"11000000000101000000000000000101",
"10111000000000000000000000000000",
"10000001000100000000000000000001",
"10100000110011000000000000000000",
"01000000000000000000001000101111",
"10111000000000000000000000000000",
"00000000100100001000000000000000",
"10000000100010000000000001000001",
"10111000000101000000000000000000",
"10111000000100000000000000000000",
"10111000000011000000000000000000",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"10000000100110000000000000000000",
"10111000000010000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"01000100000000000000001010010100",
"01000100000000000000001010000010",
"10010000000000000000000000000000",
"10000000000000000000000010010110",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001010111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000101",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010010",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"01000100000000000000001010010100",
"01000100000000000000001010000010",
"10010000000000000000000000000000",
"10000000000000000000000010010110",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001001100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000101",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001001000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"10010000000000000000000000000000",
"10000000000000000000000010011011",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100001111000000000000000000",
"10110100001110000000000000000000",
"10010011101110000000000000000000",
"10000011101110000000000000000110",
"10010011111111000000000000000000",
"11001011111110000000000000001010",
"10110011110000000000000011001000",
"10010000000000000000000011111111",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000100000",
"01000100000000000000000100101001",
"10000011111111000000000000000001",
"01000000000000000000001010000111",
"10111000001110000000000000000000",
"10111000001111000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000011010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000100000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10000111111111000000000000000001",
"10110011110000000000000011001000",
"10110100000000000000000000000000",
"10010000000000000000000011111111",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10111000000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10100100000000000000000000000000",
"10010000000000000000000011111111",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10000000010001000000000011010100",
"10110100000000000000000000000000",
"10000000010000000000000000000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10111000000000000000000000000000",
"01000100000000000000000100101001",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000111110100",
"10010000010001000000000000000000",
"11000000010000000000000000000100",
"01000100000000000000000101001010",
"10000100000000000000000000000001",
"01000000000000000000001011001010",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10110100000010000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000011010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"10010000100010000000000000000000",
"10000000100010000000000000000001",
"11001000100001000000000000000100",
"01000100000000000000000100101001",
"10000000100010000000000000000001",
"01000000000000000000001011011100",
"10111000000010000000000000000000",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000010010100",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000001001000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001000101",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001001100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000001010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000111010",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"00000000000001000001000000000000",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10110100000010000000000000000000",
"10110100000011000000000000000000",
"10110100000100000000000000000000",
"10110100000101000000000000000000",
"10110100000110000000000000000000",
"10110100000111000000000000000000",
"10110100001000000000000000000000",
"10110100001001000000000000000000",
"10110100001010000000000000000000",
"10110100001011000000000000000000",
"10110100001100000000000000000000",
"10110100001101000000000000000000",
"10110100001110000000000000000000",
"10110100001111000000000000000000",
"01000100000000000000010001100000",
"10010000010001000000000000000000",
"10010000000000000000000000000000",
"10010001010101000000000000000000",
"10000001010101000000000000010011",
"11000000010101000000000100000000",
"10000000010010000000000000000001",
"10000000010011000000000000000010",
"10000000010100000000000000000011",
"01000100000000000000010000010011",
"10000000010000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000010000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10000000100000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000010",
"01000100000000000000000100101001",
"10000000100000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10000000110000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000000110000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000101",
"01000100000000000000000100101001",
"01000100000000000000010001111110",
"01000100000000000000010010001010",
"10000000010000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000010000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10000000100000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000010",
"01000100000000000000000100101001",
"10000000100000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10000000110000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000000110000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000101",
"01000100000000000000000100101001",
"01000100000000000000010001111110",
"01000100000000000000010011100100",
"10000000010000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000010000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10000000100000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000010",
"01000100000000000000000100101001",
"10000000100000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10000000110000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000000110000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000101",
"01000100000000000000000100101001",
"01000100000000000000010001111110",
"01000100000000000000010100111110",
"10000000010000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000000010000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000000100000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000100000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10000000110000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000010",
"01000100000000000000000100101001",
"10000000110000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"01000100000000000000010001111110",
"01000100000000000000010110001111",
"10000000010000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000110",
"01000100000000000000000100101001",
"10000000010000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000110",
"01000100000000000000000100101001",
"10000000100000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000100000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10000000110000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000010",
"01000100000000000000000100101001",
"10000000110000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10000001000000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000001000000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000101",
"01000100000000000000000100101001",
"01000100000000000000010001111110",
"01000100000000000000010111111000",
"10000000100000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000100000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10000000110000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000010",
"01000100000000000000000100101001",
"10000000110000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10000001000000000000000010000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000100",
"01000100000000000000000100101001",
"10000001000000000000000011000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000101",
"01000100000000000000000100101001",
"01000100000000000000010001111110",
"10000000010001000000000000000001",
"01000000000000000000001100010010",
"10111000001111000000000000000000",
"10111000001110000000000000000000",
"10111000001101000000000000000000",
"10111000001100000000000000000000",
"10111000001011000000000000000000",
"10111000001010000000000000000000",
"10111000001001000000000000000000",
"10111000001000000000000000000000",
"10111000000111000000000000000000",
"10111000000110000000000000000000",
"10111000000101000000000000000000",
"10111000000100000000000000000000",
"10111000000011000000000000000000",
"10111000000010000000000000000000",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010100000000000000000000000100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"11010000000000000000000000000000",
"01000100000000000000000101001010",
"10000000000000000000000000111000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000001100",
"01000100000000000000000100011111",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"10000000000000000000000000000110",
"01000100000000000000000100011111",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001100100",
"10010000010001000000000000000000",
"11000000000001111111110011000011",
"10000100000000000000000000000001",
"01000000000000000000000100111000",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10110100000001000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000000010100",
"10010000010001000000000000000000",
"11000000010000000000000000000100",
"01000100000000000000000101001010",
"10000100000000000000000000000001",
"01000000000000000000010010000011",
"10111000000001000000000000000000",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10010100000000000000000000000010",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010100000000000000000000000100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"10010100000000000000000000001000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"10010100000000000000000000001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010100000000000000000000000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001000000",
"01000100000000000000000100011111",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10010100000000000000000000000010",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010100000000000000000000000100",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010100000000000000000000000001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010100000000000000000000000001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001000000",
"01000100000000000000000100011111",
"01000100000000000000000101001010",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000011",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000000111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000001111",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011111",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010100000000000000000000000001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011100",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000011110",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010100000000000000000000001000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"10000000000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"10010100000000000000000000010000",
"01000100000000000000000100101001",
"10010000000000000000000000000000",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"01000100000000000000000100101001",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000010000000000000000000",
"10010011010010000000000000000111",
"10110100000001000000000000000000",
"10001000100001000000000000000011",
"10000000010001000000000000001101",
"10000000010000000000000000000000",
"10111000000001000000000000000000",
"10111000000010000000000000000000",
"01001000000000000000000000000000",--
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10000000000000000000000011001111",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10000000000000000000000010100011",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001000001",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000","10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000010100011",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011100010",
"01000100000000000000000100010010",
"01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001111100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"10111000000000000000000000000000",
"01001000000000000000000000000000",
"10110100000110000000000000000000",
"10110100000011000000000000000000",
"10110100000010000000000000000000",
"10110100000001000000000000000000",
"10110100000101000000000000000000","10110100000101000000000000000000",
"10010000110011000000000000000000",
"10010000010001000000000000000000",
"10010100010001000000000000000001",
"00000001010001001001000000000000",
"10010011111111000000000000000000",
"11000000101111000000000000000110",
"10100101010101000000000000000000",
"10000000110011000000000000000001",
"01000000000000000000000011111000",
"01000100000000000000000100010010","01000100000000000000000100111101",
"10010000000000000000000000000000",
"10000000000000000000000001011111",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"01000100000000000000000100011100",
"10010000000000000000000000000000",
"10000000000000000000000011001111",
"01000100000000000000000100010010"
);


instruction<= ins_mem(conv_integer(unsigned(pc)));
end Behavioral;

